
module day5_tb ();

  logic clk;
  logic reset;

  logic [2:0] cnt_o;

  day5 DAY5 (.*);

  always begin
    clk = 1'b0;
    #5;
    clk = 1'b1;
    #5;
  end

  initial begin
    reset = 1'b1;
    @(posedge clk);
    @(posedge clk);
    reset = 1'b0;
    for (int i=0; i<30; i++)
      @(posedge clk);
    $finish();
  end

endmodule