module tb;
reg clk, rst, load;
reg [2:0] parallel_in;
wire serial_out;

piso dut(clk, rst, load, parallel_in, serial_out);

	always #5 clk = !clk;
 
  initial begin 
  clk=0;
  	#2;
	rst=1;
	#2;
	rst=0;
  end
    
 initial begin
    #5;
    load= 1'b1;
    parallel_in= 3'b001;
    #10 load= 1'b0;
    #30 load= 1'b1;
    parallel_in= 3'b100;
    #10 load= 1'b0;
    #30 load= 1'b1;
    parallel_in= 3'b101;
    #10 load= 1'b0;
	
	#20;
	$finish;
    end
    
endmodule